entity Hazard_Unit is
    Port (
        POPM : in std_logic;
    );
end Hazard_Unit;