entity Hazard_Unit is
    Port (
        POPM : in std_logic;
        PUSM : in std_logic;
        Mem : in std_logic;
        IsIMM : in std_logic;
        RTI:
    );
end Hazard_Unit;