entity Hazard_Unit is
    Port (
        Pop
    );
end Hazard_Unit;