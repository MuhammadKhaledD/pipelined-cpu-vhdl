entity Hazard_Unit is
    Port (
        
    );
end Hazard_Unit;