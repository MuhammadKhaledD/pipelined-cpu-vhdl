entity Ha