entity Haza